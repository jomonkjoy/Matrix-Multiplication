byte_write_spram #(
) (
);

endmodule
