module matrix_multiply #(
) (
);

endmodule
