module multiply_acc #(
) (
);

endmodule
